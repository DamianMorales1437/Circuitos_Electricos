** Profile: "SCHEMATIC1-lab5_3"  [ C:\Users\daxda\OneDrive\Documentos\Universidad\Dispositivos electronicos\laboratorios\lab5_2180389_B02\lab5_2180389_b02-pspicefiles\schematic1\lab5_3.sim ] 

** Creating circuit file "lab5_3.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../lab5_2180389_b02-pspicefiles/lab5_2180389_b02.lib" 
* From [PSPICE NETLIST] section of C:\Users\daxda\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 30m 0 0.1u 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
