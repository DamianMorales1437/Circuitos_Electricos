** Profile: "SCHEMATIC1-lab2_sumador"  [ C:\Users\Demian\Documents\universidad\dispositivos electronicos\laboratorios\lab2_2180389_B02-PSpiceFiles\SCHEMATIC1\lab2_sumador.sim ] 

** Creating circuit file "lab2_sumador.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "D:/Lite Small/tools/capture/library/pspice/nat_semi.lib" 
* From [PSPICE NETLIST] section of C:\SPB_DATA\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 3ms 0 0.1u 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
