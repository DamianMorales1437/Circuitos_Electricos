** Profile: "SCHEMATIC1-curva pasabajas"  [ C:\Users\daxda\OneDrive\Documentos\Universidad\Dispositivos electronicos\laboratorios\lab4_2180389_B02\lab4_2180389_b02-pspicefiles\schematic1\curva pasabajas.sim ] 

** Creating circuit file "curva pasabajas.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "D:/Programas/universidad/orcad/tools/capture/library/pspice/nat_semi.lib" 
* From [PSPICE NETLIST] section of C:\Users\daxda\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 100 1 1Meg
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
