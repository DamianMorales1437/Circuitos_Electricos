** Profile: "SCHEMATIC1-1"  [ C:\USERS\DAXDA\ONEDRIVE\DOCUMENTOS\UNIVERSIDAD\DISPOSITIVOS ELECTRONICOS\LABORATORIOS 2\LAB8_2180389_B04\LAB8_2180389_BO4-PSpiceFiles\SCHEMATIC1\1.sim ] 

** Creating circuit file "1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../lab8_2180389_bo4-pspicefiles/lab8_2180389_bo4.lib" 
* From [PSPICE NETLIST] section of C:\Users\daxda\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN V_V1 -24 12 0.1 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
