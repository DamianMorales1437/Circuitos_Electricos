** Profile: "SCHEMATIC1-simlab1_2"  [ C:\Users\Demian\Documents\universidad\dispositivos\laboratorios\lab1_2180389_B02\lab1-PSpiceFiles\SCHEMATIC1\simlab1_2.sim ] 

** Creating circuit file "simlab1_2.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "D:/Lite Small/tools/capture/library/pspice/opamp.lib" 
* From [PSPICE NETLIST] section of C:\SPB_DATA\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 3ms 0 10u 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
